--test bench

